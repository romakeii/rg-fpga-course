`timescale 1ns / 1ps

// Дешифратор - комбинационная схема, преобразующая
// n-разрядный код числа на входе в код разрядности 2^n
// На выходной порт, индекс которого соответствует значению на входе, выдается "1";
// на остальные выходные порты выдается "0"
// Пример схемы:
//    |‾‾‾‾‾‾‾|
//    |decoder|
//    |       |
// 1--|i0   o0|--0
//    |     o1|--1
//    |     o2|--0
// 0--|i1   o3|--0
//    |_______|

// Реализовать дешифратор с разрядностью входа, равной 2 битам
// Названия входных/выходных портов - "in"/"out"
// Использовать процедурный блок always_comb и оператор case
// Выходные значения описать двоичными литералами

module decoder_1of4 (
// Описание портов
);
// Описание логики
endmodule

// Реализовать дешифратор, размерность входной шины которого задается парамертом "IN_WIDTH"
// Названия входных/выходных портов - "in"/"out"
// Использовать процедурный блок always_comb и оператор []

module decoder_prm #(
// Описание параметров
) (
// Описание портов
);
// Описание логики
endmodule

// Неполный дешифратор - дешифратор, имеющий n разрядов на входе
// и меньше, чем 2^n разрядов на выходе
// Т.е. это такой дешифратор, у которого НЕ ДЛЯ ВСЕХ возможных входных значений
// существует выход с соответствующим индексом

// Реализовать дешифратор, размерность ВЫходной шины которого задается параметром "OUT_WIDTH"
// Размерность входной шины должна выражаться через параметр OUT_WIDTH при помощи системной функции $clog2()
// Названия входных/выходных портов - "in"/"out"
// Использовать процедурный блок always_comb и оператор []
// Предусмотреть случай использования модуля в качестве неполного дешифратора (например, когда при инстанцировании задали OUT_WIDTH = 3):
// в этом случае при установке значения на входе, не имеющего соответствующего выхода, все выходы дешифратора должны устанавливаться в 0

module decoder_oprm #(
// Описание параметров
) (
// Описание портов
);
// Описание логики
endmodule
