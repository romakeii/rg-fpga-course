`timescale 1ns / 1ns

// Реализовать тестбенч для проверки модуля srl_bus
// Сформировать тактовый сигнал, сброс и входное воздействие для тестируемого модуля
// Реализовать проверку ожидаемого результата на выходе тестируемого модуля
// При реализации формирования входного воздействия и проверки использовать код из модуля srl_bit_tb, поместив
// этот код в task в файл tasks.sv и подключив его к данному файлу
// В коде модуля srl_bus_tb использовать вызов этого task

module srl_bus_tb;

endmodule

// Переписать код модуля srl_bit_tb с использованием task из файла tasks.sv
