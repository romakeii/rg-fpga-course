`timescale 1ns / 1ps

// Дешифратор - комбинационная схема, преобразующая
// n-разрядный код числа на входе в код разрядности 2^n
// На выходной порт, индекс которого соответствует значению на входе, выдается "1";
// на остальные выходные порты выдается "0"
// Пример схемы:
//    |‾‾‾‾‾‾‾|
//    |decoder|
//    |       |
// 1--|i0   o0|--0
//    |     o1|--1
//    |     o2|--0
// 0--|i1   o3|--0
//    |_______|

// Реализовать дешифратор с разрядностью входа, равной 2 битам
// Названия входных/выходных портов - "in"/"out"
// Использовать процедурный блок always_comb и оператор case
// Выходные значения описать двоичными литералами

module decoder_1of4 (

// Описание портов
    input  logic [1 : 0] in,
    output logic [3 : 0] out

);

// Описание логики
    always_comb begin
        case (in)
            2'b00   : out = 4'b0001;
            2'b01   : out = 4'b0010;
            2'b10   : out = 4'b0100;
            2'b11   : out = 4'b1000;
            default : out = 4'b0000;
        endcase
    end

endmodule

// Реализовать дешифратор, размерность входной шины которого задается парамертом "IN_WIDTH"
// Названия входных/выходных портов - "in"/"out"
// Использовать процедурный блок always_comb и оператор []

module decoder_prm #(

// Описание параметров
    parameter IN_WIDTH = 2

) (

// Описание портов
    input logic [IN_WIDTH - 1 : 0] in,
    output logic [2**IN_WIDTH - 1 : 0] out

);

// Описание логики
    always_comb begin
        out = '0; // необязательная строка, т.к. следующей строкой исчерпывающе описываются все выходные значения при любых возможных входах;
        // это происходит потому, что параметром задается размер входной шины, а размер выходной вычисляется исходя из его значения,
        // т.е. не может быть такого значения на входе, которое не соответствует какому-то из индексов выходной шины
        out[in] = 1'b1;
    end

endmodule

// Неполный дешифратор - дешифратор, имеющий n разрядов на входе
// и меньше, чем 2^n разрядов на выходе
// Т.е. это такой дешифратор, у которого НЕ ДЛЯ ВСЕХ возможных входных значений
// существует выход с соответствующим индексом

// Реализовать дешифратор, размерность ВЫходной шины которого задается параметром "OUT_WIDTH"
// Размерность входной шины должна выражаться через параметр OUT_WIDTH при помощи системной функции $clog2()
// Названия входных/выходных портов - "in"/"out"
// Использовать процедурный блок always_comb и оператор []
// Предусмотреть случай использования модуля в качестве неполного дешифратора (например, когда при инстанцировании задали OUT_WIDTH = 3):
// в этом случае при установке значения на входе, не имеющего соответствующего выхода, все выходы дешифратора должны устанавливаться в 0

module decoder_oprm #(

// Описание параметров
    parameter OUT_WIDTH = 4
) (

// Описание портов
    input logic [$clog2(OUT_WIDTH) - 1 : 0] in,
    output logic [OUT_WIDTH - 1 : 0] out
);

// Описание логики
    always_comb begin
        out = '0; // в отличие от дешифратора decoder_prm, в описании данного модуля эту строку писать обязательно, чтобы не получить защелку при синтезе;
        // в данном модуле параметром задается размер выходной шины, а размер входной вычисляется исходя из его значения,
        // т.е., в зависимости от значения параметра, могут существовать такие значения на входе, которое не соответствует ни одному из индексов выходной шины
        // Следовательно, опиав выходы ТОЛЬКО с использованием строки ниже, мы можем (если зададим параметр != степени 2) не учесть некоторые варианты входного значения
        // и не определим выход для такого значения
        out[in] = 1'b1;
    end

endmodule
