`timescale 1ns / 1ns

task automatic make_in (

);

endtask

task compare (

);

endtask
