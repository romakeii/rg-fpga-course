`timescale 1ns / 1ps

// Реализовать линию задержки однобитового сигнала
// Длина линии задержки (количество тактов задержки) должна задаваться параметром
// Требуемые порты:
// входы клока, синхронного сброса и данных (1 бит),
// выход данных (1 бит)

// Shift register line (SRL)
module srl_bit #(
// Описание параметров
) (
// Описание портов
);
// Описание логики
endmodule
