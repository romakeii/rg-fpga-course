`timescale 1ns / 1ps

// Реализовать устройство логического сдвига, размерности входной и выходной шин которого задаются параметром "WIDTH"
// Сигнал "in" - входная шина, "out" - выходная шина, "drc" - выбор направления сдвига (0 - вправо, 1 - влево)
// Количество разрядов сдвига должно задаваться параметром "SHIFT"
// Использовать непрерывное присваивание с оператором "?:" (для выбора направления сдвига) и операторы логического сдвига (>> и <<)

module shift_operator #(
    parameter   WIDTH = 16,
    parameter   SHIFT = 1
) (
    input logic     [WIDTH-1:0] in,
    input logic                 drc,
    output logic    [WIDTH-1:0] out
);
    assign out = drc ? (in << SHIFT) : (in >> SHIFT);

endmodule

// Реализовать устройство логического сдвига, размерности входной и выходной шин которого задаются параметром "WIDTH"
// Сигнал "in" - входная шина, "out" - выходная шина, "drc" - выбор направления сдвига (0 - вправо, 1 - влево)
// Количество разрядов сдвига должно задаваться параметром "SHIFT"
// Использовать непрерывное присваивание с оператором "?:" (для выбора направления сдвига) и оператор конкатенации {}

module shift_with_concat #(
    parameter   WIDTH = 16,
    parameter   SHIFT = 1
) (
    input logic     [WIDTH-1:0] in,
    input logic                 drc,
    output logic    [WIDTH-1:0] out
);

    // Внутри оператора конкатенации слева у шины "in" обозначать диапазон индексов не обязательно,
    // т.к. старшая часть, не помещающаяся в разрядную сетку шины "out", будет отброшена автоматически
    // Внутри оператора конкатенации справа диапазон индексов шины "in" нужно указывать явно,
    // т.к. в этом случае должна быть отброшена МЛАДШАЯ часть
    assign out = drc ? {in, {SHIFT{1'b0}}} : {{SHIFT{1'b0}}, in[WIDTH - 1 : SHIFT]};

endmodule
