`timescale 1ns / 1ns

// Реализовать тестбенч для проверки модуля srl_bit
// Сформировать тактовый сигнал, сброс и входное воздействие для тестируемого модуля
// Реализовать проверку ожидаемого результата на выходе тестируемого модуля

module srl_bit_tb;
// Описание логики
endmodule

// Выполнить задание из файла srl_bus.sv
