`timescale 1ns / 1ps

// Реализовать устройство логического сдвига, размерности входной и выходной шин которого задаются параметром "WIDTH"
// Сигнал "in" - входная шина, "out" - выходная шина, "drc" - выбор направления сдвига (0 - вправо, 1 - влево)
// Количество разрядов сдвига должно задаваться параметром "SHIFT"
// Использовать непрерывное присваивание с оператором "?:" (для выбора направления сдвига) и операторы логического сдвига (>> и <<)

module shift_operator #(
// Описание параметров
) (
// Описание портов
);
// Описание логики
endmodule

// Реализовать устройство логического сдвига, размерности входной и выходной шин которого задаются параметром "WIDTH"
// Сигнал "in" - входная шина, "out" - выходная шина, "drc" - выбор направления сдвига (0 - вправо, 1 - влево)
// Количество разрядов сдвига должно задаваться параметром "SHIFT"
// Использовать непрерывное присваивание с оператором "?:" (для выбора направления сдвига) и оператор конкатенации {}

module shift_with_concat #(
// Описание параметров
) (
// Описание портов
);
// Описание логики
endmodule
