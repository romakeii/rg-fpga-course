`timescale 1ns / 1ps

// Реализовать линию задержки для шины
// Длина линии задержки (количество тактов задержки) должна задаваться параметром
// Ширина шины должна задаваться параметром
// Требуемые порты:
// входы клока, синхронного сброса и данных (количество бит задается параметром),
// выход данных (количество бит задается параметром)
// Для реализации использовать generage блок и инстанцированный модуль srl_bit
// из файла srl_bit.sv

module srl_bus #(
// Описание параметров
) (
// Описание портов
);
// Описание логики
endmodule
